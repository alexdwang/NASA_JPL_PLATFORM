Title: AD590 / Pre Rad / T= 300.15K = 27C
*

*Voltage Source
VIN 1 0 DC 0V

*Umbrella circuit
X1 1 2 AD590_sc
ROUT 2 0 1m

*Input
.dc VIN 0 30 0.01

*Output
.print dc format=noindex file=AD590_Prerad_27C_V1.txt
+ V(1)
+ I(ROUT)

*Subcircuit
.subckt AD590_sc IN OUT

*Capacitance: C<name> <+ node> <- node> [model name] <value> + [IC=<initial value>]
c1 1 8 26p

*Resistance: R<name> <+ node> <- node> [model name] <value>
r1 IN 4 260
r2 IN 3 1040
r3 5 16 5000
r4 11 5 11000
r5 12 OUT 146
r6 15 OUT 820

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q11 1 5 12 QNMOD 35 temp=27
Q10 5 5 12 QNMOD 35 temp=27
Q9 6 5 15 QNMOD 280 temp=27
Q6 7 7 IN QLPMOD 10 temp=27
Q4 1 8 4 QLPMOD 10 temp=27
Q3 1 8 4 QLPMOD 10 temp=27
Q5 8 8 3 QLPMOD 10 temp=27
Q2 6 8 4 QLPMOD 10 temp=27
Q1 6 8 4 QLPMOD 10 temp=27
Q7 7 6 11 QNMOD 10 temp=27
Q8 8 1 11 QNMOD 10 temp=27

*JFET: J<name> <drain> <gate> <source> <model name> [area value]
J1 8 16 11 NJF_TYP

*end of the subcircuit
.ends

*Library
* npn prerad off ctp 3b
.model QNMOD NPN (
+ IS = 1.68208E-16
+ BF = 84.058    NF = 0.986787 VAF = 351.9861415
+ IKF = 9.86E-3  NK = 0.47574  ISE = 7.1029E-15
+ NE = 2.06453   BR = 0.697    NR = 2
+ VAR = 100      IKR = 0.1     ISC = 1E-17
+ NC = 2         RB = 140.86   IRB = 1E-3
+ RBM = 50       RE = 2        RC = 250.75)

*lpnp prerad off ctp 3b
.model QLPMOD PNP (
+ IS = 8.70964E-16
+ BF = 786.9		NF = 0.99                           VAF = 36.3423711
+ IKF = 6.30957E-5       NK = 0.52                           ISE = 9.54993E-17
+ NE = 1.27089           BR = 0.697                          NR = 2
+ VAR = 100              IKR = 0.1                           ISC = 1E-17
+ NC = 2                 RB = 758.578                        IRB = 3.6E-5
+ RBM = 100              RE = 4.096                           RC = 1)

*JFET
.model NJF_TYP NJF (
+ VTO = -1.0	BETA = 6.2E-4	LAMBDA = 0.003
+ RD = 0.01      RS = 1e-4
+ CGS = 3E-12    CGD=1.5E-12     IS=5E-10)

*end of the netlist
.end
