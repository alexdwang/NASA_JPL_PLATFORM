Title: LT1175 / Line Regulation / ABM / 2.5krad / T= 300.15K = 27C

*Input Voltage Source
V2 4 0 DC 0V

*Schematic name: LT1175 core
****************************
*Subcircuit
*X1 VCC VEE VREF
X1 0 4 5 BG_sc

*X4 V+ V- VCC VEE VO
X4 6 5 0 4 7 OPAMP_sc

*Resistance: R<name> <+ node> <- node> [model name] <value>
r1 0 6 350k
r2 6 1 100k
rLIM 3 4 0.001

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q1 1 2 3 QNMOD 1000
Q2 0 7 2 QNMOD 10

*Parameters
***********
*PRE_RAD
.PARAM a1=-39.30421
.PARAM b1=48.21879
.PARAM c1=-15.6477

*2.5krad
.PARAM a2=-39.12298
.PARAM b2=53.5479
.PARAM c2=-21.84106

*SCALE
.PARAM scale1=1
.PARAM scale2=1
.PARAM scale3=1
.PARAM scale4=0.1

.PARAM scale6=20
.PARAM scale7=20
.PARAM scale8=1
.PARAM scale9=10
.PARAM scale10=10

*Function
*********
*DeltaIb = 1*(exp(a2+(b2*Veb)+(c2*(Veb*Veb))) - exp(a1+(b1*Veb)+(c1*(Veb*Veb))))
*.func deltaIb(x) {scale*(exp(a2+(b2*x)+(c2*(pow(x,2)))) - exp(a1+(b1*x)+(c1*(pow(x,2)))))}
.func deltaIb1(x) {scale1*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb2(x) {scale2*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb3(x) {scale3*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb4(x) {scale4*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}

.func deltaIb6(x) {scale6*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb7(x) {scale7*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb8(x) {scale8*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb9(x) {scale9*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}
.func deltaIb10(x) {scale10*(exp(a2+(b2*x)+(c2*(x*x))) - exp(a1+(b1*x)+(c1*(x*x))))}

*Input
.dc V2 0 -20 -0.1

*Output
.print dc format=noindex file=LT1175_Prerad_LineRegulation_V12_ABM_2krad.txt
+ V(4)
+ V(1)


*Schematic name: BG_sc
**********************
.subckt BG_sc VCC VEE VREF
*Voltage Controlled Current Source BG
B1 VCC 2 I={deltaIb1(V(VCC)-V(2))}
B2 1 2 I={deltaIb2(V(1)-V(2))}
B3 9 5 I={deltaIb3(V(9)-V(5))}
B4 8 5 I={deltaIb4(V(8)-V(5))}

*Resistance: R<name> <+ node> <- node> [model name] <value>
r1 VCC 1 10k
r2 1 8 2.93e6
r3 8 9 109k
r4 4 VEE 600
r5 6 VEE 600

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q1 2 2 VCC QLPMOD 1
Q2 3 2 1 QLPMOD 1
Q3 12 5 9 QLPMOD 1
Q4 11 5 8 QLPMOD 0.1
Q5 12 12 7 QNMOD 1
Q6 11 12 7 QNMOD 1
Q7 VCC 5 7 QNMOD 1
Q8 3 3 4 QNMOD 1
Q9 7 3 6 QNMOD 1

*Voltage Controlled Voltage Source: E<name> <+ node> <-node> <+ controlling node> <- controlling node> <gain>
E1 VCC VREF VCC 5 1

*Independent Current Source: I<name> <+ node> <-node> [[DC] <value>]
I1 2 0 DC 3.23uA

*end of the BG_sc subcircuit
.ends BG_sc


*Schematic name: OPAMP_sc
*************************
.subckt OPAMP_sc V10 V11 VCC VEE VO

*Voltage Controlled Current Source OPAMP
B6 5 V10 I={deltaIb6(V(5)-V(V10))}
B7 5 V11 I={deltaIb7(V(5)-V(V11))}
B8 6 VCC I={deltaIb8(V(6)-V(VCC))}
B9 6 VCC I={deltaIb9(V(6)-V(VCC))}
B10 6 VCC I={deltaIb10(V(6)-V(VCC))}

*Resistance: R<name> <+ node> <- node> [model name] <value>
r1 7 VEE 4.7k
r2 3 VEE 4.7k
r3 VO VEE 60k
r4 11 VEE 60k

*Capacitance: C<name> <+ node> <- node> [model name] <value> + [IC=<initial value>]
C1 1 9 0.0056p

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q1 1 11 VEE QNMOD 10
Q2 VCC 1 VO QNMOD 1
Q3 VCC 9 11 QNMOD 1
Q4 9 4 7 QNMOD 1
Q5 4 4 3 QNMOD 1
Q6 9 V10 5 QLPMOD 20
Q7 4 V11 5 QLPMOD 20
Q8 6 6 VCC QLPMOD 1
Q9 5 6 VCC QLPMOD 10
Q10 1 6 VCC QLPMOD 10

*Independent Current Source: I<name> <+ node> <-node> [[DC] <value>]
I1 6 0 DC 1.4u

*end of the OPAMP_sc subcircuit
.ends OPAMP_sc

*Library
********
* npn prerad off ctp 3b
.model QNMOD NPN (              
+ IS = 1.68208E-16
+ BF = 84.058    NF = 0.986787 VAF = 351.9861415
+ IKF = 9.86E-3  NK = 0.47574  ISE = 7.1029E-15
+ NE = 2.06453   BR = 0.697    NR = 2
+ VAR = 100      IKR = 0.1     ISC = 1E-17
+ NC = 2         RB = 140.86   IRB = 1E-3
+ RBM = 50       RE = 2        RC = 250.75)

*lpnp prerad off ctp 3b
.model QLPMOD PNP (             
+ IS = 8.70964E-16
+ BF = 786.9		NF = 0.99                           VAF = 36.3423711
+ IKF = 6.30957E-5       NK = 0.52                           ISE = 9.54993E-17
+ NE = 1.27089           BR = 0.697                          NR = 2
+ VAR = 100              IKR = 0.1                           ISC = 1E-17
+ NC = 2                 RB = 758.578                        IRB = 3.6E-5
+ RBM = 100              RE = 4.096                           RC = 1)

*end of the netlist
.end
