Title: AD590 / 20k / Current source / T= 300.15K = 27C
*************************************

*Input voltage source
***************
VIN 2 0 DC 0V

*Circuit Core
*************
XZ 2 20 AD590
R0 20 0 1m

*Parameters
***********
*PRE_RAD_PNP
.PARAM a1=-41.935
.PARAM b1=47.6314
.PARAM c1=-11.045

*20krad_PNP
.PARAM a2=-32.249
.PARAM b2=35.6571
.PARAM c2=-9.1636

*PRE_RAD_NPN
.PARAM a3=-39.91
.PARAM b3=40.6194
.PARAM c3=-4.4288

*20krad_NPN
.PARAM a4=-34.92
.PARAM b4=30.4499
.PARAM c4=1.11115

*SCALE
.PARAM scale1=10
.PARAM scale2=10
.PARAM scale3=10
.PARAM scale4=10
.PARAM scale5=10
.PARAM scale6=10
.PARAM scale7=10
.PARAM scale8=10
.PARAM scale9=280
.PARAM scale10=35
.PARAM scale11=35

*Function
*********
*DeltaIb = 1*(exp(a2+(b2*Veb)+(c2*(Veb*Veb))) - exp(a1+(b1*Veb)+(c1*(Veb*Veb))))
*.func deltaIb(x) {scale*(exp(a2+(b2*x)+(c2*(pow(x,2)))) - exp(a1+(b1*x)+(c1*(pow(x,2)))))}
*PNP
.func deltaIb1(x) {scale1*((exp(a2+(b2*x)+(c2*(x*x)))) - (exp(a1+(b1*x)+(c1*(x*x)))))}
.func deltaIb2(x) {scale2*((exp(a2+(b2*x)+(c2*(x*x)))) - (exp(a1+(b1*x)+(c1*(x*x)))))}
.func deltaIb3(x) {scale3*((exp(a2+(b2*x)+(c2*(x*x)))) - (exp(a1+(b1*x)+(c1*(x*x)))))}
.func deltaIb4(x) {scale4*((exp(a2+(b2*x)+(c2*(x*x)))) - (exp(a1+(b1*x)+(c1*(x*x)))))}
.func deltaIb5(x) {scale5*((exp(a2+(b2*x)+(c2*(x*x)))) - (exp(a1+(b1*x)+(c1*(x*x)))))}
.func deltaIb6(x) {scale6*((exp(a2+(b2*x)+(c2*(x*x)))) - (exp(a1+(b1*x)+(c1*(x*x)))))}

*NPN
.func deltaIb7(x) {scale7*((exp(a4+(b4*x)+(c4*(x*x)))) - (exp(a3+(b3*x)+(c3*(x*x)))))}
.func deltaIb8(x) {scale8*((exp(a4+(b4*x)+(c4*(x*x)))) - (exp(a3+(b3*x)+(c3*(x*x)))))}
.func deltaIb9(x) {scale9*((exp(a4+(b4*x)+(c4*(x*x)))) - (exp(a3+(b3*x)+(c3*(x*x)))))}
.func deltaIb10(x) {scale10*((exp(a4+(b4*x)+(c4*(x*x)))) - (exp(a3+(b3*x)+(c3*(x*x)))))}
.func deltaIb11(x) {scale11*((exp(a4+(b4*x)+(c4*(x*x)))) - (exp(a3+(b3*x)+(c3*(x*x)))))}

*Input
******
.dc VIN 0 30 0.01

*Output
*******
.print dc format=noindex file=AD590_27C_20k_CurrentSource.txt
+ V(2)
+ I(R0)

*Subcircuit
************
.subckt AD590 2 20

*Voltage Controlled Current Source
*PNP
B1 4 8 I={deltaIb1(V(4)-V(8))}
B2 4 8 I={deltaIb2(V(4)-V(8))}
B3 4 8 I={deltaIb3(V(4)-V(8))}
B4 4 8 I={deltaIb4(V(4)-V(8))}
B5 3 8 I={deltaIb5(V(3)-V(8))}
B6 2 7 I={deltaIb6(V(2)-V(7))}
*NPN
B7 6 11 I={deltaIb7(V(6,11))}
B8 1 11 I={deltaIb8(V(1,11))}
B9 5 15 I={deltaIb9(V(5,15))}
B10 5 12 I={deltaIb10(V(5,12))}
B11 5 12 I={deltaIb11(V(5,12))}

*Capacitance: C<name> <+ node> <- node> [model name] <value> + [IC=<initial value>]
c1 1 8 26p

*Resistance: R<name> <+ node> <- node> [model name] <value>
r1 2 4 260
r2 2 3 1040
r3 5 16 5000
r4 11 5 11000
r5 12 20 146
r6 15 20 820

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q11 1 5 12 QNMOD 35 temp=27
Q10 5 5 12 QNMOD 35 temp=27
Q9 6 5 15 QNMOD 280 temp=27
Q6 7 7 2 QLPMOD 10 temp=27
Q4 1 8 4 QLPMOD 10 temp=27
Q3 1 8 4 QLPMOD 10 temp=27
Q5 8 8 3 QLPMOD 10 temp=27
Q2 6 8 4 QLPMOD 10 temp=27
Q1 6 8 4 QLPMOD 10 temp=27
Q7 7 6 11 QNMOD 10 temp=27
Q8 8 1 11 QNMOD 10 temp=27

*JFET: J<name> <drain> <gate> <source> <model name> [area value]
J1 8 16 11 NJF_TYP

*end of the subcircuit 
.ends

*Library
********
* npn prerad off ctp 3b
.model QNMOD NPN (              
+ IS = 1.68208E-16
+ BF = 84.058    NF = 0.986787 VAF = 351.9861415
+ IKF = 9.86E-3  NK = 0.47574  ISE = 7.1029E-15
+ NE = 2.06453   BR = 0.697    NR = 2
+ VAR = 100      IKR = 0.1     ISC = 1E-17
+ NC = 2         RB = 140.86   IRB = 1E-3
+ RBM = 50       RE = 2        RC = 250.75)

*lpnp prerad off ctp 3b
.model QLPMOD PNP (             
+ IS = 8.70964E-16
+ BF = 786.9		NF = 0.99                           VAF = 36.3423711
+ IKF = 6.30957E-5       NK = 0.52                           ISE = 9.54993E-17
+ NE = 1.27089           BR = 0.697                          NR = 2
+ VAR = 100              IKR = 0.1                           ISC = 1E-17
+ NC = 2                 RB = 758.578                        IRB = 3.6E-5
+ RBM = 100              RE = 4.096                           RC = 1) 

*JFET
.model NJF_TYP NJF (
+ VTO = -1.0	BETA = 6.2E-4	LAMBDA = 0.003 
+ RD = 0.01      RS = 1e-4 
+ CGS = 3E-12    CGD=1.5E-12     IS=5E-10)

*end of the netlist
.end
